`include "Mux_4X1.v"
`timescale 1ns/1ps

module Mux_4X1_TB;
 reg i0,i1,i2,i3;
 reg s0,s1;
 wire Y;

 Mux_4X1 DUT (i0,i1,i2,i3,s0,s1,Y);

 initial begin
   $monitor("TIME = %0dns  i0 = %0d   i1 = %0d   i2 = %0d   i3 = %0d   s0 = %0d   s1 = %0d   Y = %0d",$time,i0,i1,i2,i3,s0,s1,Y);

        i0 = 0; i1 = 0; i2 = 0; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 0; s0 = 1; s1 = 1;

	 
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 0; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 0; i2 = 1; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 0; i2 = 1; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 0; i2 = 1; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 1; i2 = 0; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 1; i2 = 0; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 0; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 1; i2 = 1; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 0; i1 = 1; i2 = 1; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 0; i1 = 1; i2 = 1; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 0; i2 = 0; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 0; i2 = 0; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 0; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 0; i2 = 1; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 0; i2 = 1; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 0; i2 = 1; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 1; i2 = 0; i3 = 0; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 0; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 0; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 0; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 1; i2 = 0; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 0; i3 = 1; s0 = 1; s1 = 1;


#10     i0 = 1; i1 = 1; i2 = 1; i3 = 1; s0 = 0; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 1; i3 = 1; s0 = 0; s1 = 1;
#10     i0 = 1; i1 = 1; i2 = 1; i3 = 1; s0 = 1; s1 = 0;
#10     i0 = 1; i1 = 1; i2 = 1; i3 = 1; s0 = 1; s1 = 1;

#10;
$finish;
end
endmodule
